module seven_seg_decoder(
	[3:0] in,
	[7:0] seg);
	
	input in;
	output seg;
	
	
endmodule